`timescale 1ns / 1ps

package uart_pkg;

  typedef enum {
    NONE,
    EVEN,
    ODD
  } parity_t;

endpackage
